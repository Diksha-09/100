`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

// 
//////////////////////////////////////////////////////////////////////////////////


module MUX_4X1(S, I, Y);
    input [1:0]S;
    input[3:0] I;
    output Y;
    reg Y;
    always @(*)
    begin
    if (S[0] == 0 && S[1] == 0)
    Y <= I[0];
    if (S[1] == 0 && S[0] == 1)
    Y <= I[1];
    if (S[0] == 0 && S[1] == 1)
    Y <= I[2];
    if (S[0] == 1 && S[1] == 1)
    Y <= I[3];
    end
    endmodule
